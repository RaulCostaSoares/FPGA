module Calculadora(
    input logic [3:0] cmd,  // comando: dígito ou operador
    input logic reset,
    input logic clock, 

    output logic [1:0] status, // estado atual
    output logic [3:0] pos,     // posição do display 
    output logic [3:0] dig      // dígito para o display
);

    typedef enum logic [1:0] {ERRO, PRONTA, OCUPADA} statetype;
    statetype estados;

    reg [31:0] reg1, reg2, saida, contador;
    reg [3:0] op;
    reg set_op, flag, flag_div;
    reg [3:0] pos_atual; // contador de posição de dígito

    assign status = estados; 

    always @(posedge clock) begin
        if (reset) begin
            estados  <= PRONTA;
            op       <= 4'b1010;
            dig      <= 0;
            pos      <= 0;
            set_op   <= 0;
            flag     <= 0;
            flag_div <= 0;
            reg1     <= 0;
            reg2     <= 0;
            saida    <= 0;
            contador <= 0;
            pos_atual <= 0;
        end else begin
            case (estados)
                PRONTA: begin
                    if (cmd < 10 && !set_op) begin
                        reg1 <= (reg1 * 10) + cmd;
                        dig <= cmd;
                        pos <= pos; // mantém posição atual (ou pode incrementar se quiser)
                        flag <= 1;
                    end 
                    else if (cmd < 10 && set_op) begin 
                        reg2 <= (reg2 * 10) + cmd;
                        dig <= cmd;
                        pos <= pos; 
                        flag <= 1;
                    end 
                    else if (cmd == 4'b1110) begin
                        case (op)
                            4'b1010: begin
                                saida <= reg1 + reg2;
                                estados <= OCUPADA;
                                pos_atual <= 0;
                            end                
                            4'b1011: begin
                                saida <= reg1 - reg2;
                                estados <= OCUPADA;
                                pos_atual <= 0;
                            end  
                            4'b1100: begin
                                if (reg1 == 0 || reg2 == 0) begin
                                    estados <= ERRO;
                                end else begin
                                    saida <= 0;
                                    contador <= 0;
                                    estados <= OCUPADA;
                                    pos_atual <= 0;
                                end
                            end
                            default: estados <= PRONTA;
                        endcase
                    end 
                    else if ((!set_op && reg1 > 32'd99999999) || (set_op && reg2 > 32'd99999999)) begin
                        estados <= ERRO;
                        pos <= 0;
                    end 
                    else begin
                        op <= cmd;
                        set_op <= 1;
                    end
                end

                ERRO: begin
                    if (cmd == 4'b1111) begin
                        estados  <= PRONTA;
                        reg1     <= 0;
                        reg2     <= 0;
                        saida    <= 0;
                        op       <= 0;
                        set_op   <= 0;
                        contador <= 0;
                        dig      <= 0;
                        pos      <= 0;
                        pos_atual <= 0;
                    end
                end

                OCUPADA: begin
                    if (op == 4'b1100 && contador < reg2) begin
                        saida <= saida + reg1;
                        contador <= contador + 1;
                    end 
                    else begin
                        if (saida > 32'd99999999) begin
                            estados <= ERRO;
                        end 
                        else begin
                            case (pos_atual)
                                0: dig <= (saida / 10000000) % 10;
                                1: dig <= (saida / 1000000) % 10;
                                2: dig <= (saida / 100000) % 10;
                                3: dig <= (saida / 10000) % 10;
                                4: dig <= (saida / 1000) % 10;
                                5: dig <= (saida / 100) % 10;
                                6: dig <= (saida / 10) % 10;
                                7: dig <= saida % 10;
                                default: dig <= 0;
                            endcase
                            
                            pos <= pos_atual;
                            pos_atual <= pos_atual + 1;

                            if (pos_atual == 8) begin
                                estados <= PRONTA;
                                reg1 <= 0;
                                reg2 <= 0;
                                saida <= 0;
                                op <= 4'b1010;
                                set_op <= 0;
                                contador <= 0;
                                pos_atual <= 0;
                            end
                        end
                    end
                end

            endcase
        end
    end

endmodule
